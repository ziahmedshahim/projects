module barrel_shifter_8bit_tb;
  reg [7:0] in;
  reg [2:0] ctrl;
  wire [7:0] out; 
  
barrel_shifter_8bit uut(.in(in), .ctrl(ctrl), .out(out));
  
initial 
 begin
    $display($time, " << Starting the Simulation >>");
        in= 8'd0;  ctrl=3'd0; //no shift
    #10 in=8'b10000000; ctrl= 3'd4; //shift 4 bit
    #10 in=8'b10000000; ctrl= 3'd2; //shift 2 bit
    #10 in=8'b10000000; ctrl= 3'd1; //shift by 1 bit
    #10 in=8'b10000000; ctrl= 3'd7; //shift by 7bit
  end
    initial begin
      $monitor("Input=%d, Control=%d, Output=%b",in,ctrl,out);
    end
    initial begin
    $dumpfile("waveform.vcd");
    $dumpvars();
    end
endmodule
